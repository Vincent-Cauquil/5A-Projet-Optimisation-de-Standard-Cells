* XOR2 Energy
.title XOR2 Energy

.lib /path/to/sky130.lib.spice tt

.param SUPPLY=1.8
.param TEMP=27
.param CLOAD=10f
.param FREQ=100MEG

.temp {TEMP}

VVDD VDD 0 DC {SUPPLY}
VVSS VSS 0 DC 0

CL Y 0 {CLOAD}

X1 A B Y VDD VSS sky130_fd_sc_hd__xor2_1

* Signaux à FREQ
VA A 0 PULSE(0 {SUPPLY} 0 100p 100p {1/(2*FREQ)} {1/FREQ})
VB B 0 PULSE(0 {SUPPLY} 0 100p 100p {1/(4*FREQ)} {1/(2*FREQ)})

.tran 1p {10/FREQ}

* Mesures sur les dernières périodes (stable)
.meas tran Iavg_total AVG i(VVDD) FROM={8/FREQ} TO={10/FREQ}
.meas tran Pavg_total PARAM='{-Iavg_total*SUPPLY}'
.meas tran Etot_avg PARAM='{Pavg_total/FREQ}'

.control
run
quit
.endc

.end