* Caractérisation de l'énergie totale - XOR2_1
* PDK Sky130 - Bibliothèque sky130_fd_sc_hd

.lib "~/.ciel/sky130/libs.tech/ngspice/sky130.lib.spice" tt
.include "~/.ciel/sky130/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

*======================================================================
* Paramètres de simulation
*======================================================================
.param SUPPLY = 1.8
.param TEMP = 27
.temp TEMP

* Paramètres de timing
.param trise = 100p
.param tfall = 100p
.param tpulse = 5n

*======================================================================
* Sources d'alimentation
*======================================================================
Vdd vdd 0 dc SUPPLY
Vss vss 0 dc 0

*======================================================================
* Cellule sous test
*======================================================================
Xxor2 A B Y vdd vss sky130_fd_sc_hd__xor2_1

*======================================================================
* Charge de sortie
*======================================================================
Cload Y 0 10f

*======================================================================
* Stimuli - Séquence optimale (même que délai)
*======================================================================

.param t0 = 1n
.param t1 = 't0+tpulse'
.param t2 = 't1+tpulse'
.param t3 = 't2+tpulse'
.param t4 = 't3+tpulse'
.param tend = 't4+tpulse'

* Signal A
VA A 0 PWL(
+ 0 0
+ t0 0
+ t1 0
+ 't1+trise' 0
+ t2 0
+ 't2+trise' SUPPLY
+ t3 SUPPLY
+ t4 SUPPLY
+ 't4+tfall' 0
+ tend 0
+ )

* Signal B
VB B 0 PWL(
+ 0 0
+ t0 0
+ t1 0
+ 't1+trise' SUPPLY
+ t2 SUPPLY
+ t3 SUPPLY
+ 't3+tfall' 0
+ t4 0
+ tend 0
+ )

*======================================================================
* Mesures d'énergie totale (selon formule (6) du document)
* Etotal = ∫ [P_VDD(t) + P_VA(t) + P_VB(t)] dt
*======================================================================

* Transition t1: B↗⇒Y↗ (A=0, état 00→01)
.measure tran t1_start param='t1'
.measure tran t1_end param='t1+1n'
.measure tran E_vdd_t1 INTEG '-I(Vdd)*SUPPLY' FROM='t1_start' TO='t1_end'
.measure tran E_vA_t1 INTEG '-I(VA)*0' FROM='t1_start' TO='t1_end'
.measure tran E_vB_t1 INTEG '-I(VB)*SUPPLY' FROM='t1_start' TO='t1_end'
.measure tran E_total_t1 param='E_vdd_t1+E_vA_t1+E_vB_t1'

* Transition t2: A↗⇒Y↘ (B=1, état 01→11)
.measure tran t2_start param='t2'
.measure tran t2_end param='t2+1n'
.measure tran E_vdd_t2 INTEG '-I(Vdd)*SUPPLY' FROM='t2_start' TO='t2_end'
.measure tran E_vA_t2 INTEG '-I(VA)*SUPPLY' FROM='t2_start' TO='t2_end'
.measure tran E_vB_t2 INTEG '-I(VB)*SUPPLY' FROM='t2_start' TO='t2_end'
.measure tran E_total_t2 param='E_vdd_t2+E_vA_t2+E_vB_t2'

* Transition t3: B↘⇒Y↗ (A=1, état 11→10)
.measure tran t3_start param='t3'
.measure tran t3_end param='t3+1n'
.measure tran E_vdd_t3 INTEG '-I(Vdd)*SUPPLY' FROM='t3_start' TO='t3_end'
.measure tran E_vA_t3 INTEG '-I(VA)*SUPPLY' FROM='t3_start' TO='t3_end'
.measure tran E_vB_t3 INTEG '-I(VB)*0' FROM='t3_start' TO='t3_end'
.measure tran E_total_t3 param='E_vdd_t3+E_vA_t3+E_vB_t3'

* Transition t4: A↘⇒Y↘ (B=0, état 10→00)
.measure tran t4_start param='t4'
.measure tran t4_end param='t4+1n'
.measure tran E_vdd_t4 INTEG '-I(Vdd)*SUPPLY' FROM='t4_start' TO='t4_end'
.measure tran E_vA_t4 INTEG '-I(VA)*0' FROM='t4_start' TO='t4_end'
.measure tran E_vB_t4 INTEG '-I(VB)*0' FROM='t4_start' TO='t4_end'
.measure tran E_total_t4 param='E_vdd_t4+E_vA_t4+E_vB_t4'

* Énergie totale moyenne par transition
.measure tran E_avg param='(E_total_t1+E_total_t2+E_total_t3+E_total_t4)/4'

*======================================================================
* Simulation
*======================================================================
.tran 10p 'tend'

.control
run
plot v(A)+4 v(B)+2 v(Y)
plot -I(Vdd)
print E_total_t1 E_total_t2 E_total_t3 E_total_t4 E_avg
.endc

.end
