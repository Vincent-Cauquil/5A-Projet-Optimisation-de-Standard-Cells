* Caractérisation de la consommation statique - XOR2_1
* PDK Sky130 - Bibliothèque sky130_fd_sc_hd

.lib "~/.ciel/sky130/libs.tech/ngspice/sky130.lib.spice" tt
.include "~/.ciel/sky130/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

*======================================================================
* Paramètres de simulation
*======================================================================
.param SUPPLY = 1.8
.param TEMP = 27
.temp TEMP

* Temps de stabilisation
.param tstab = 10n
.param tduration = 5n

*======================================================================
* Sources d'alimentation
*======================================================================
Vdd vdd 0 dc SUPPLY
Vss vss 0 dc 0

*======================================================================
* Cellule sous test
*======================================================================
Xxor2 A B Y vdd vss sky130_fd_sc_hd__xor2_1

*======================================================================
* Pas de charge nécessaire pour consommation statique
*======================================================================

*======================================================================
* Stimuli - Tous les états
* État 1: A=0 B=0 Y=0
* État 2: A=0 B=1 Y=1
* État 3: A=1 B=0 Y=1
* État 4: A=1 B=1 Y=0
*======================================================================

.param t1 = tstab
.param t2 = 't1+tduration'
.param t3 = 't2+tduration'
.param t4 = 't3+tduration'
.param tend = 't4+tduration'

* Signal A
VA A 0 PWL(
+ 0 0
+ t1 0
+ t2 0
+ t3 SUPPLY
+ t4 SUPPLY
+ tend SUPPLY
+ )

* Signal B
VB B 0 PWL(
+ 0 0
+ t1 0
+ t2 SUPPLY
+ t3 0
+ t4 SUPPLY
+ tend SUPPLY
+ )

*======================================================================
* Mesures de consommation statique (selon formule (5) du document)
* L(A,B) = P(VDD) + P(VA) + P(VB)
* L(A,B) = -VDD*I(VDD) - VA*I(VA) - VB*I(VB)
*======================================================================

* État 1: A=0, B=0
.measure tran I_vdd_00 AVG I(Vdd) FROM='t1' TO='t2'
.measure tran I_vA_00 AVG I(VA) FROM='t1' TO='t2'
.measure tran I_vB_00 AVG I(VB) FROM='t1' TO='t2'
.measure tran L_00 param='-SUPPLY*I_vdd_00 - 0*I_vA_00 - 0*I_vB_00'

* État 2: A=0, B=1
.measure tran I_vdd_01 AVG I(Vdd) FROM='t2' TO='t3'
.measure tran I_vA_01 AVG I(VA) FROM='t2' TO='t3'
.measure tran I_vB_01 AVG I(VB) FROM='t2' TO='t3'
.measure tran L_01 param='-SUPPLY*I_vdd_01 - 0*I_vA_01 - SUPPLY*I_vB_01'

* État 3: A=1, B=0
.measure tran I_vdd_10 AVG I(Vdd) FROM='t3' TO='t4'
.measure tran I_vA_10 AVG I(VA) FROM='t3' TO='t4'
.measure tran I_vB_10 AVG I(VB) FROM='t3' TO='t4'
.measure tran L_10 param='-SUPPLY*I_vdd_10 - SUPPLY*I_vA_10 - 0*I_vB_10'

* État 4: A=1, B=1
.measure tran I_vdd_11 AVG I(Vdd) FROM='t4' TO='tend'
.measure tran I_vA_11 AVG I(VA) FROM='t4' TO='tend'
.measure tran I_vB_11 AVG I(VB) FROM='t4' TO='tend'
.measure tran L_11 param='-SUPPLY*I_vdd_11 - SUPPLY*I_vA_11 - SUPPLY*I_vB_11'

* Consommation statique moyenne
.measure tran L_avg param='(L_00+L_01+L_10+L_11)/4'

*======================================================================
* Simulation
*======================================================================
.tran 10p 'tend'

.control
run
plot v(A)+4 v(B)+2 v(Y)
plot I(Vdd)
print L_00 L_01 L_10 L_11 L_avg
.endc

.end
