* Caractérisation de la consommation dynamique - XOR2_1
* PDK Sky130 - Bibliothèque sky130_fd_sc_hd
* Cette netlist mesure aussi la consommation statique (selon l'énoncé)

.lib "~/.ciel/sky130/libs.tech/ngspice/sky130.lib.spice" tt
.include "~/.ciel/sky130/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

*======================================================================
* Paramètres de simulation
*======================================================================
.param SUPPLY = 1.8
.param TEMP = 27
.temp TEMP

* Paramètres de timing
.param trise = 100p
.param tfall = 100p
.param tstab = 10n
.param tduration = 5n
.param tpulse = 5n

*======================================================================
* Sources d'alimentation
*======================================================================
Vdd vdd 0 dc SUPPLY
Vss vss 0 dc 0

*======================================================================
* Cellule sous test
*======================================================================
Xxor2 A B Y vdd vss sky130_fd_sc_hd__xor2_1

*======================================================================
* Charge de sortie
*======================================================================
Cload Y 0 10f

*======================================================================
* PHASE 1: Mesure consommation statique (tous les états)
* PHASE 2: Mesure énergie totale (transitions)
*======================================================================

* Phase 1: États statiques
.param t1_static = tstab
.param t2_static = 't1_static+tduration'
.param t3_static = 't2_static+tduration'
.param t4_static = 't3_static+tduration'

* Phase 2: Transitions dynamiques
.param t_dyn_start = 't4_static+tduration'
.param t1_dyn = 't_dyn_start'
.param t2_dyn = 't1_dyn+tpulse'
.param t3_dyn = 't2_dyn+tpulse'
.param t4_dyn = 't3_dyn+tpulse'
.param tend = 't4_dyn+tpulse'

*======================================================================
* Stimuli
*======================================================================

* Signal A
VA A 0 PWL(
+ 0 0
+ t1_static 0
+ t2_static 0
+ t3_static SUPPLY
+ t4_static SUPPLY
+ t_dyn_start 0
+ t1_dyn 0
+ t2_dyn 0
+ 't2_dyn+trise' SUPPLY
+ t3_dyn SUPPLY
+ t4_dyn SUPPLY
+ 't4_dyn+tfall' 0
+ tend 0
+ )

* Signal B
VB B 0 PWL(
+ 0 0
+ t1_static 0
+ t2_static SUPPLY
+ t3_static 0
+ t4_static SUPPLY
+ t_dyn_start 0
+ t1_dyn 0
+ 't1_dyn+trise' SUPPLY
+ t2_dyn SUPPLY
+ t3_dyn SUPPLY
+ 't3_dyn+tfall' 0
+ t4_dyn 0
+ tend 0
+ )

*======================================================================
* MESURES PHASE 1: Consommation statique (formule (5))
*======================================================================

* État 1: A=0, B=0
.measure tran I_vdd_00 AVG I(Vdd) FROM='t1_static' TO='t2_static'
.measure tran I_vA_00 AVG I(VA) FROM='t1_static' TO='t2_static'
.measure tran I_vB_00 AVG I(VB) FROM='t1_static' TO='t2_static'
.measure tran L_00 param='-SUPPLY*I_vdd_00 - 0*I_vA_00 - 0*I_vB_00'

* État 2: A=0, B=1
.measure tran I_vdd_01 AVG I(Vdd) FROM='t2_static' TO='t3_static'
.measure tran I_vA_01 AVG I(VA) FROM='t2_static' TO='t3_static'
.measure tran I_vB_01 AVG I(VB) FROM='t2_static' TO='t3_static'
.measure tran L_01 param='-SUPPLY*I_vdd_01 - 0*I_vA_01 - SUPPLY*I_vB_01'

* État 3: A=1, B=0
.measure tran I_vdd_10 AVG I(Vdd) FROM='t3_static' TO='t4_static'
.measure tran I_vA_10 AVG I(VA) FROM='t3_static' TO='t4_static'
.measure tran I_vB_10 AVG I(VB) FROM='t3_static' TO='t4_static'
.measure tran L_10 param='-SUPPLY*I_vdd_10 - SUPPLY*I_vA_10 - 0*I_vB_10'

* État 4: A=1, B=1
.measure tran I_vdd_11 AVG I(Vdd) FROM='t4_static' TO='t_dyn_start'
.measure tran I_vA_11 AVG I(VA) FROM='t4_static' TO='t_dyn_start'
.measure tran I_vB_11 AVG I(VB) FROM='t4_static' TO='t_dyn_start'
.measure tran L_11 param='-SUPPLY*I_vdd_11 - SUPPLY*I_vA_11 - SUPPLY*I_vB_11'

*======================================================================
* MESURES PHASE 2: Énergie totale (formule (6))
*======================================================================

* Transition t1: état 00→01 (B↗⇒Y↗)
.measure tran t1_start param='t1_dyn'
.measure tran t1_end param='t1_dyn+1n'
.measure tran E_total_t1 INTEG '-I(Vdd)*SUPPLY-I(VA)*0-I(VB)*SUPPLY' FROM='t1_start' TO='t1_end'

* Transition t2: état 01→11 (A↗⇒Y↘)
.measure tran t2_start param='t2_dyn'
.measure tran t2_end param='t2_dyn+1n'
.measure tran E_total_t2 INTEG '-I(Vdd)*SUPPLY-I(VA)*SUPPLY-I(VB)*SUPPLY' FROM='t2_start' TO='t2_end'

* Transition t3: état 11→10 (B↘⇒Y↗)
.measure tran t3_start param='t3_dyn'
.measure tran t3_end param='t3_dyn+1n'
.measure tran E_total_t3 INTEG '-I(Vdd)*SUPPLY-I(VA)*SUPPLY-I(VB)*0' FROM='t3_start' TO='t3_end'

* Transition t4: état 10→00 (A↘⇒Y↘)
.measure tran t4_start param='t4_dyn'
.measure tran t4_end param='t4_dyn+1n'
.measure tran E_total_t4 INTEG '-I(Vdd)*SUPPLY-I(VA)*0-I(VB)*0' FROM='t4_start' TO='t4_end'

*======================================================================
* Calcul consommation dynamique (formule (7))
* Edyn = Etotal - L(S0)×(t1-t0) - L(S1)×(t2-t1)
*======================================================================

* Transition 1: 00→01
.measure tran dt1 param='1n'
.measure tran E_static_t1_before param='L_00*dt1'
.measure tran E_static_t1_after param='L_01*0'
.measure tran Edyn_t1 param='E_total_t1-E_static_t1_before-E_static_t1_after'

* Transition 2: 01→11
.measure tran dt2 param='1n'
.measure tran E_static_t2_before param='L_01*dt2'
.measure tran E_static_t2_after param='L_11*0'
.measure tran Edyn_t2 param='E_total_t2-E_static_t2_before-E_static_t2_after'

* Transition 3: 11→10
.measure tran dt3 param='1n'
.measure tran E_static_t3_before param='L_11*dt3'
.measure tran E_static_t3_after param='L_10*0'
.measure tran Edyn_t3 param='E_total_t3-E_static_t3_before-E_static_t3_after'

* Transition 4: 10→00
.measure tran dt4 param='1n'
.measure tran E_static_t4_before param='L_10*dt4'
.measure tran E_static_t4_after param='L_00*0'
.measure tran Edyn_t4 param='E_total_t4-E_static_t4_before-E_static_t4_after'

* Énergie dynamique moyenne
.measure tran Edyn_avg param='(Edyn_t1+Edyn_t2+Edyn_t3+Edyn_t4)/4'

*======================================================================
* Simulation
*======================================================================
.tran 10p 'tend'

.control
run
plot v(A)+4 v(B)+2 v(Y)
plot -I(Vdd)
echo "=== CONSOMMATION STATIQUE ==="
print L_00 L_01 L_10 L_11
echo "=== ÉNERGIE TOTALE ==="
print E_total_t1 E_total_t2 E_total_t3 E_total_t4
echo "=== CONSOMMATION DYNAMIQUE ==="
print Edyn_t1 Edyn_t2 Edyn_t3 Edyn_t4 Edyn_avg
.endc

.end
